/*
This is a Moore state machine with two states, one input, and one output. Implement this state machine. Notice that the reset state is B.

This exercise is the same as fsm1, but using synchronous reset.
*/

// Note the Verilog-1995 module declaration syntax here:
module top_module(clk, reset, in, out);
    input clk;
    input reset;    // Synchronous reset to state B
    input in;
    output out;		//  
    reg out;

    parameter A=1'b0, B=1'b1;		// Fill in state name declarations
    reg present_state, next_state;

    always @(posedge clk) begin
        if (reset) begin  
            present_state = B;		// Fill in reset logic
        end else begin
            case (present_state)
                A: next_state = in ? A : B;
                B: next_state = in ? B : A;		// Fill in state transition logic
            endcase

            // State flip-flops
            present_state = next_state;   
        end
            case (present_state)
                A: out = 1'b0;		// Fill in output logic
                B: out = 1'b1;
            endcase
    end

endmodule
